library verilog;
use verilog.vl_types.all;
entity sum_product is
end sum_product;
