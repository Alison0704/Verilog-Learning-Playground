library verilog;
use verilog.vl_types.all;
entity hello_world is
end hello_world;
